module main

fn test_solve_a() {
	input := ['1,9,10,3,2,3,11,0,99,30,40,50']
	assert solve_a(input, -1, -1) == 3500
}

// Not possible to test solve_b() without actual test data
// which I'm not gonna make public...
// Feel free to PR
