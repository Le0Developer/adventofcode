module main

fn test_solve_a() {
	inputs := ['2 * 3 + (4 * 5)', '5 + (8 * 3 + 9 + 3 * 4 * 3)', '5 * 9 * (7 * 3 * 3 + 9 * 3 + (8 + 6 * 4))',
		'((2 + 4 * 9) * (6 + 9 * 8 + 6) + 6) + 2 + 4 * 2',
	]
	assert solve_a(inputs) == 26335
}

fn test_solve_b() {
	inputs := ['2 * 3 + (4 * 5)', '5 + (8 * 3 + 9 + 3 * 4 * 3)', '5 * 9 * (7 * 3 * 3 + 9 * 3 + (8 + 6 * 4))',
		'((2 + 4 * 9) * (6 + 9 * 8 + 6) + 6) + 2 + 4 * 2',
	]
	assert solve_b(inputs) == 693891
}
