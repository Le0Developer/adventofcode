module main

fn test_solve_a() {
	input := ['100000-250000']
	assert solve_a(input) == 1877
}

fn test_solve_b() {
	input := ['100000-250000']
	assert solve_b(input) == 1374
}
