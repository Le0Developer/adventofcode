module main

fn test_solve_a() {
	inputs := ['12', '14', '1969', '100756']
	assert solve_a(inputs) == 34241
}

fn test_solve_b() {
	inputs := ['12', '14', '1969', '100756']
	assert solve_b(inputs) == 51316
}
