module main

import flag
import os

fn challenge_a(input_lines []string) ?i64 {
	mut previous := input_lines[0].int()
	mut total := 0
	for line in input_lines {
		as_int := line.int()
		if as_int > previous {
			total++
		}
		previous = as_int
	}
	return total
}

fn challenge_b(input_lines []string) ?i64 {
	mut previous1 := input_lines[0].int()
	mut previous2 := input_lines[1].int()
	mut previous_sum := input_lines[0].int() + input_lines[1].int() + input_lines[2].int()
	mut total := 0
	for line in input_lines[2..] {
		as_int := line.int()
		sum := previous1 + previous2 + as_int
		if sum > previous_sum {
			total++
		}
		previous_sum = sum
		previous1 = previous2
		previous2 = as_int
	}
	return total
}

fn main() {
	mut fp := flag.new_flag_parser(os.args)
	fp.application('AdventOfCode 202_ day __')
	fp.version('v0.1.0')
	fp.skip_executable()
	fp.limit_free_args_to_exactly(1) ?
	is_b := fp.bool('b', `b`, false, 'b challenge')
	// more options here
	additional_args := fp.finalize() or {
		eprintln(err)
		println(fp.usage())
		return
	}
	input_filename := additional_args[0]
	input_lines := os.read_lines(input_filename) ?
	solution := if !is_b { challenge_a(input_lines) ? } else { challenge_b(input_lines) ? }
	println('Solution is $solution')
}
