module main

fn test_solve_a() {
	inputs := [16, 10, 15, 5, 1, 11, 7, 19, 6, 12, 4]
	assert solve_a(inputs) == 35
}

fn test_solve_b() {
	inputs := [16, 10, 15, 5, 1, 11, 7, 19, 6, 12, 4]
	assert solve_b(inputs) == 8
}
